* SKY130 1.8V NMOS wrapper
* Wraps sky130_fd_pr__nfet_01v8 with simplified interface
* Dimensions in um (with NGspice scale=1e-6)

.subckt nfet_01v8 d g s b
.param w=1 l=0.15 nf=1 mult=1
XM d g s b sky130_fd_pr__nfet_01v8 w={w} l={l} nf={nf} mult={mult}
.ends nfet_01v8

* SKY130 MiM Capacitor wrapper (M4-M5)
* Wraps sky130_fd_pr__cap_mim_m3_2 with simplified interface
* Requires: .lib sky130.lib.spice tt

.subckt cap_mim_m4 PLUS MINUS
.param w=10 l=10 mult=1
XC PLUS MINUS sky130_fd_pr__cap_mim_m3_2 w={w} l={l} mult={mult}
.ends cap_mim_m4
